
module INSTRUCTION_FETCH(
	clk,
	rst,
	jump,
	branch,
	jump_addr,
	branch_addr,

	PC,
	IR
);

input clk, rst, jump, branch;
input [31:0] jump_addr, branch_addr;

output reg 	[31:0] PC;
output reg 	[31:0] IR;

reg [31:0] instruction [127:0];
//output instruction
always @(posedge clk or posedge rst)
begin
	if(rst) begin
		IR <= 32'd0;
		instruction[ 0] = 32'b100011_00000_00010_00000_00000_000000;//lw $2 imm($s0)  = $S2 <= mem[imm + S0]
        instruction[ 1] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[ 2] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[ 3] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[ 4] = 32'b000000_00010_00000_00101_00000_100000;    //add(add $5, $2, $0)
        instruction[ 5] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[ 6] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[ 7] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)        
    
        instruction[ 8] = 32'b000000_00000_00001_00100_00000_100000;    //add(add $4, $0, $1)
        instruction[ 9] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[10] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[11] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        //comp_b
        instruction[12] = 32'b000000_00000_00001_00100_00000_100000;    //add(add $4, $0, $1)
        instruction[13] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[14] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[15] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
    
        instruction[16] = 32'b000000_00101_00001_00101_00000_100000;    //add(add $5, $5, $1)
        instruction[17] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[18] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[19] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
//        $display("DONE");
        instruction[20] = 32'b000000_00101_00000_00011_00000_100000;    //add(add $3, $0, $5)
        instruction[21] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[22] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[23] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        //adiv
        instruction[24] = 32'b000000_00100_00001_00100_00000_100000;    //add(add $4, $4, $1)
        instruction[25] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[26] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[27] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[28] = 32'b000000_00101_00000_00011_00000_100000;    //add(add $3, $5, $0)
        instruction[29] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[30] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[31] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        //judgeP
        instruction[32] = 32'b000000_00011_00100_00011_00000_100010;    //sub(sub $3, $3, $4)
        instruction[33] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[34] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[35] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[36] = 32'b000000_00100_00011_00110_00000_101010;    //slt(slt $6, $4, $3)
        instruction[37] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[38] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[39] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[40] = 32'b000101_00110_00000_11111_11111_110111;    //bne(bne $6, $0, judgeP)
        instruction[41] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[42] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[43] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        //checkB
        instruction[44] = 32'b000100_00011_00100_11111_11111_011111;    //beq(beq $3, $4, comp_b)
        instruction[45] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[46] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[47] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[48] = 32'b000101_00101_00100_11111_11111_100011;    //bne(bne $4, $5, adiv)
        instruction[49] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[50] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[51] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        //printB
        instruction[52] = 32'b101011_00000_00101_00000_00000_000010;    //sw $3 imm($s2) = mem[imm + S2] <= $3
        instruction[53] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[54] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[55] = 32'b000000_00000_00000_00000_00000_100000; //NOP
    
        instruction[56] = 32'b000000_00010_00000_00101_00000_100000;    //add(add $5, $2, $0)
        instruction[57] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[58] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[59] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[60] = 32'b000000_00000_00001_00100_00000_100000;    //add(add $4, $0, $1)
        instruction[61] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[62] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[63] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
    
        
        
        //comp_s
        instruction[64] = 32'b000000_00000_00001_00100_00000_100000;    //add(add $4, $0, $1)
        instruction[65] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[66] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[67] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[68] = 32'b000000_00101_00001_00101_00000_100010;    //sub(sub $5, $5, $1)
        instruction[69] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[70] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[71] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[72] = 32'b000000_00101_00000_00011_00000_100000;    //add(add $3, $0, $5)
        instruction[73] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[74] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[75] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        //adiv_s
        instruction[76] = 32'b000000_00100_00001_00100_00000_100000;    //add(add $4, $4, $1)
        instruction[77] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[78] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[79] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[80] = 32'b000000_00101_00000_00011_00000_100000;    //add(add $3, $5, $0)
        instruction[81] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[82] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[83] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        //judgePs
        instruction[84] = 32'b000000_00011_00100_00011_00000_100010;    //sub(sub $3, $3, $4)
        instruction[85] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[86] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[87] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[88] = 32'b000000_00100_00011_00110_00000_101010;    //slt(slt $6, $4, $3)
        instruction[89] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[90] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[91] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
    
        instruction[92] = 32'b000101_00110_00000_11111_11111_110111;    //bne(bne $6, $0, judgePs)
        instruction[93] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[94] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[95] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        //check
        instruction[96] = 32'b000100_00011_00100_11111_11111_011111;    //beq(beq $3, $4, comp_s)
        instruction[97] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[98] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[99] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        
        instruction[100] = 32'b000101_00101_00100_11111_11111_100011;    //bne(bne $4, $5, adiv)
        instruction[101] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[102] = 32'b000000_00000_00000_00000_00000_100000;//NOP(add $0, $0, $0)
        instruction[103] = 32'b000000_00000_00000_00000_00000_100000;//NOP(add $0, $0, $0)
        //printS
        instruction[104] = 32'b101011_00000_00101_00000_00000_000011;    //sw $5 imm($s2) = mem[imm + S2] <= $5
        instruction[105] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[106] = 32'b000000_00000_00000_00000_00000_100000;    //NOP(add $0, $0, $0)
        instruction[107] = 32'b000000_00000_00000_00000_00000_100000; //NOP
        
	end
	else begin
		if(PC[10:2]<=8'd127) 
		  IR <= instruction[PC[10:2]]; //(0, 4, 8, ...) => (0, 1, 2, ...)
		//else
		  //IR <= IR;
	end
end

// output program counter
always @(posedge clk or posedge rst)
begin
	if(rst)
		PC <= 32'd0;
	else begin
	   if(PC[10:2]<8'd127) 
	       PC <= (branch) ? branch_addr : ( (jump) ? jump_addr : (PC+4)) ;
	   //else
	       //PC <= PC;
	end
end

endmodule